* C:\Users\telep\Documents\Documents\ECL\1A\UEs\STI\tc0\Elec\2_NMOS_AMP\AMP.sch

* Schematics Version 9.1 - Web Update 1
* Sun Jan 21 10:44:42 2018



** Analysis setup **
.tran 1us 10ms 0 1us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "C:\Program Files\OrCAD_Demo\PSpice\Library\eea.lib"
.lib "nom.lib"

.INC "AMP.net"
.INC "AMP.als"


.probe


.END
