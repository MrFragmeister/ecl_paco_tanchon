* C:\Users\telep\Documents\Documents\ECL\1A\UEs\STI\tc0\Elec\7_NE555_astab\NE555_Astable.sch

* Schematics Version 9.1 - Web Update 1
* Sun Jan 21 15:56:59 2018



** Analysis setup **
.tran 1ns 50us 0 1ns
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "C:\Program Files\OrCAD_Demo\PSpice\Library\eea.lib"
.lib "nom.lib"

.INC "NE555_Astable.net"
.INC "NE555_Astable.als"


.probe


.END
