* C:\Users\telep\Documents\Documents\ECL\1A\UEs\STI\tc0\Elec\Circuits\TD5\Adder_BCD_Student.sch

* Schematics Version 9.1 - Web Update 1
* Mon Jan 22 09:04:42 2018



** Analysis setup **
.tran 0ns 400us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "C:\Program Files\OrCAD_Demo\PSpice\Library\eea.lib"
.lib "nom.lib"

.INC "Adder_BCD_Student.net"
.INC "Adder_BCD_Student.als"


.probe


.END
