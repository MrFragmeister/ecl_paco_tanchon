* C:\Users\telep\Documents\Documents\ECL\1A\UEs\STI\tc0\Elec\5_CMOS\CMOS.sch

* Schematics Version 9.1 - Web Update 1
* Sun Jan 21 15:34:45 2018



** Analysis setup **
.DC LIN V_VIN 0 2.5 0.01 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "C:\Program Files\OrCAD_Demo\PSpice\Library\eea.lib"
.lib "nom.lib"

.INC "CMOS.net"
.INC "CMOS.als"


.probe


.END
